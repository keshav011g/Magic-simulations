magic
tech scmos
timestamp 1731217574
<< nwell >>
rect -19 -8 48 88
<< ntransistor >>
rect 60 24 62 48
rect 85 24 87 48
<< ptransistor >>
rect 1 -1 3 71
rect 27 -1 29 71
<< ndiffusion >>
rect 55 47 60 48
rect 59 25 60 47
rect 55 24 60 25
rect 62 47 67 48
rect 62 25 63 47
rect 80 46 85 48
rect 62 24 67 25
rect 84 26 85 46
rect 80 24 85 26
rect 87 46 92 48
rect 87 26 88 46
rect 87 24 92 26
<< pdiffusion >>
rect -4 63 1 71
rect 0 3 1 63
rect -4 -1 1 3
rect 3 63 8 71
rect 3 3 4 63
rect 22 64 27 71
rect 3 -1 8 3
rect 26 4 27 64
rect 22 -1 27 4
rect 29 64 34 71
rect 29 4 30 64
rect 29 -1 34 4
<< ndcontact >>
rect 55 25 59 47
rect 63 25 67 47
rect 80 26 84 46
rect 88 26 92 46
<< pdcontact >>
rect -4 3 0 63
rect 4 3 8 63
rect 22 4 26 64
rect 30 4 34 64
<< psubstratepcontact >>
rect 71 32 76 39
rect 88 13 92 18
<< nsubstratencontact >>
rect 1 79 9 84
rect 13 45 18 55
rect 13 30 18 40
rect 13 13 18 23
<< polysilicon >>
rect 1 71 3 74
rect 27 71 29 74
rect 60 48 62 51
rect 85 48 87 51
rect 60 21 62 24
rect 85 21 87 24
rect 1 -4 3 -1
rect 27 -4 29 -1
<< metal1 >>
rect -4 84 0 88
rect -4 79 1 84
rect 9 79 12 84
rect -4 63 0 79
rect 8 55 22 58
rect 8 45 13 55
rect 18 45 22 55
rect 8 40 22 45
rect 8 30 13 40
rect 18 30 22 40
rect 8 23 22 30
rect 8 13 13 23
rect 18 13 22 23
rect 8 10 22 13
rect 34 31 55 40
rect 67 39 80 46
rect 67 32 71 39
rect 76 32 80 39
rect 67 26 80 32
rect 88 18 92 26
<< labels >>
rlabel polysilicon 27 72 29 74 1 Vb2
rlabel polysilicon 60 50 62 51 1 vb3
rlabel polysilicon 85 50 87 51 1 vin
rlabel metal1 88 18 92 19 7 gnd
rlabel metal1 49 31 52 40 1 vout
rlabel metal1 -4 86 0 88 5 vdd
rlabel polysilicon 1 74 3 74 1 vb1
<< end >>
